-- NCO_tb.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity NCO_tb is
	port (
		nco_ii_0_clk_clk     : in  std_logic                     := '0';             -- nco_ii_0_clk.clk
		nco_ii_0_in_valid    : in  std_logic                     := '0';             --  nco_ii_0_in.valid
		nco_ii_0_in_data     : in  std_logic_vector(15 downto 0) := (others => '0'); --             .data
		nco_ii_0_out_data    : out std_logic_vector(23 downto 0);                    -- nco_ii_0_out.data
		nco_ii_0_out_valid   : out std_logic;                                        --             .valid
		nco_ii_0_rst_reset_n : in  std_logic                     := '0'              -- nco_ii_0_rst.reset_n
	);
end entity NCO_tb;

architecture rtl of NCO_tb is
	component NCO_tb_nco_ii_0 is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset_n   : in  std_logic                     := 'X';             -- reset_n
			clken     : in  std_logic                     := 'X';             -- valid
			phi_inc_i : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			fsin_o    : out std_logic_vector(23 downto 0);                    -- data
			out_valid : out std_logic                                         -- valid
		);
	end component NCO_tb_nco_ii_0;

	signal nco_ii_0_fsin_o : std_logic_vector(23 downto 0); -- port fragment

begin

	nco_ii_0 : component NCO_tb_nco_ii_0
		port map (
			clk                    => nco_ii_0_clk_clk,              -- clk.clk
			reset_n                => nco_ii_0_rst_reset_n,          -- rst.reset_n
			clken                  => nco_ii_0_in_valid,             --  in.valid
			phi_inc_i(15 downto 0) => nco_ii_0_in_data(15 downto 0), --    .data
			fsin_o(23 downto 0)    => nco_ii_0_fsin_o(23 downto 0),  -- out.data
			out_valid              => nco_ii_0_out_valid             --    .valid
		);

	nco_ii_0_out_data <= nco_ii_0_fsin_o(23 downto 0);

end architecture rtl; -- of NCO_tb
