-- NCO_tb.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use std.env.finish;

entity FIR_Filter_tb is
end entity FIR_Filter_tb;

architecture rtl of FIR_Filter_tb is
	component NCO_tb_nco_ii_0 is
		port (
			clk       : in  std_logic;             -- clk
			reset_n   : in  std_logic;             -- reset_n
			clken     : in  std_logic;             -- valid
			phi_inc_i : in  std_logic_vector(15 downto 0); 					  -- data
			fsin_o    : out std_logic_vector(23 downto 0);                    -- data
			out_valid : out std_logic                                         -- valid
		);
	end component NCO_tb_nco_ii_0;

	constant clk_period : time := 20 ns;
	signal clk,reset_n,valid_nco : std_logic;
	signal nco_ii_0_fsin_o : std_logic_vector(23 downto 0); -- port fragment
	signal freq_count : integer range 1 to 2**16; 
	signal Time_counter : integer range 1 to 2**16; 

begin

	clk_process :process
	begin
		 clk <= '0';
		 wait for clk_period/2;  --for 0.5 ns signal is '0'.
		 clk <= '1';
		 wait for clk_period/2;  --for next 0.5 ns signal is '1'.
	end process;

	reset_n <= '0', '1' after clk_period * 3 ;

	tb1 : process(clk)
    begin
		if reset_n = '0' then 
			freq_count <= 1;
			Time_counter <= 1;
		elsif rising_edge(clk) then 
			if freq_count = 2**16 then
				--report "Finish";
			else
				if Time_counter = 2**16/freq_count then 
					freq_count <= freq_count + 1;
					Time_counter <= 1;
				else
					Time_counter <= Time_counter + 1;
				end if;
				
			end if;
		end if;
	end process;

	SEQUENCER_PROC : process
	begin
	 
	  -- Replace this line with your testbench logic
		wait until freq_count = 2**16/2;
		report "Calling 'finish'";
		--finish;
	
	end process;

	nco_ii_0 : component NCO_tb_nco_ii_0
		port map (
			clk                    => clk,              -- clk.clk
			reset_n                => reset_n,          -- rst.reset_n
			clken                  => '1',             --  in.valid
			phi_inc_i(15 downto 0) => (others => '1'), --    .data
			fsin_o(23 downto 0)    => nco_ii_0_fsin_o(23 downto 0),  -- out.data
			out_valid              => valid_nco             --    .valid
		);


end architecture rtl; -- of NCO_tb
